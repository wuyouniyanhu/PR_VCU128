// black box definition for module_count
module count(
   input        rst,
   input        clk,
   output [3:0] count_out);
endmodule
